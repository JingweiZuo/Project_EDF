library verilog;
use verilog.vl_types.all;
entity can_bsp is
    generic(
        tp              : integer := 1
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        sample_point    : in     vl_logic;
        sampled_bit     : in     vl_logic;
        sampled_bit_q   : in     vl_logic;
        tx_point        : in     vl_logic;
        hard_sync       : in     vl_logic;
        addr            : in     vl_logic_vector(7 downto 0);
        data_in         : in     vl_logic_vector(7 downto 0);
        data_out        : out    vl_logic_vector(7 downto 0);
        fifo_selected   : in     vl_logic;
        reset_mode      : in     vl_logic;
        listen_only_mode: in     vl_logic;
        acceptance_filter_mode: in     vl_logic;
        self_test_mode  : in     vl_logic;
        release_buffer  : in     vl_logic;
        tx_request      : in     vl_logic;
        abort_tx        : in     vl_logic;
        self_rx_request : in     vl_logic;
        single_shot_transmission: in     vl_logic;
        read_arbitration_lost_capture_reg: in     vl_logic;
        read_error_code_capture_reg: in     vl_logic;
        error_capture_code: out    vl_logic_vector(7 downto 0);
        error_warning_limit: in     vl_logic_vector(7 downto 0);
        we_rx_err_cnt   : in     vl_logic;
        we_tx_err_cnt   : in     vl_logic;
        extended_mode   : in     vl_logic;
        rx_idle         : out    vl_logic;
        transmitting    : out    vl_logic;
        last_bit_of_inter: out    vl_logic;
        set_reset_mode  : out    vl_logic;
        node_bus_off    : out    vl_logic;
        error_status    : out    vl_logic;
        rx_err_cnt      : out    vl_logic_vector(8 downto 0);
        tx_err_cnt      : out    vl_logic_vector(8 downto 0);
        transmit_status : out    vl_logic;
        receive_status  : out    vl_logic;
        tx_successful   : out    vl_logic;
        need_to_tx      : out    vl_logic;
        overrun         : out    vl_logic;
        info_empty      : out    vl_logic;
        set_bus_error_irq: out    vl_logic;
        set_arbitration_lost_irq: out    vl_logic;
        arbitration_lost_capture: out    vl_logic_vector(4 downto 0);
        node_error_passive: out    vl_logic;
        node_error_active: out    vl_logic;
        rx_message_counter: out    vl_logic_vector(6 downto 0);
        acceptance_code_0: in     vl_logic_vector(7 downto 0);
        acceptance_mask_0: in     vl_logic_vector(7 downto 0);
        acceptance_code_1: in     vl_logic_vector(7 downto 0);
        acceptance_code_2: in     vl_logic_vector(7 downto 0);
        acceptance_code_3: in     vl_logic_vector(7 downto 0);
        acceptance_mask_1: in     vl_logic_vector(7 downto 0);
        acceptance_mask_2: in     vl_logic_vector(7 downto 0);
        acceptance_mask_3: in     vl_logic_vector(7 downto 0);
        tx_data_0       : in     vl_logic_vector(7 downto 0);
        tx_data_1       : in     vl_logic_vector(7 downto 0);
        tx_data_2       : in     vl_logic_vector(7 downto 0);
        tx_data_3       : in     vl_logic_vector(7 downto 0);
        tx_data_4       : in     vl_logic_vector(7 downto 0);
        tx_data_5       : in     vl_logic_vector(7 downto 0);
        tx_data_6       : in     vl_logic_vector(7 downto 0);
        tx_data_7       : in     vl_logic_vector(7 downto 0);
        tx_data_8       : in     vl_logic_vector(7 downto 0);
        tx_data_9       : in     vl_logic_vector(7 downto 0);
        tx_data_10      : in     vl_logic_vector(7 downto 0);
        tx_data_11      : in     vl_logic_vector(7 downto 0);
        tx_data_12      : in     vl_logic_vector(7 downto 0);
        tx              : out    vl_logic;
        tx_oen          : out    vl_logic
    );
end can_bsp;
