library verilog;
use verilog.vl_types.all;
entity can_registers is
    generic(
        tp              : integer := 1
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        cs              : in     vl_logic;
        we              : in     vl_logic;
        addr            : in     vl_logic_vector(7 downto 0);
        data_in         : in     vl_logic_vector(7 downto 0);
        data_out        : out    vl_logic_vector(7 downto 0);
        irq             : out    vl_logic;
        sample_point    : in     vl_logic;
        transmitting    : in     vl_logic;
        set_reset_mode  : in     vl_logic;
        node_bus_off    : in     vl_logic;
        error_status    : in     vl_logic;
        rx_err_cnt      : in     vl_logic_vector(7 downto 0);
        tx_err_cnt      : in     vl_logic_vector(7 downto 0);
        transmit_status : in     vl_logic;
        receive_status  : in     vl_logic;
        tx_successful   : in     vl_logic;
        need_to_tx      : in     vl_logic;
        overrun         : in     vl_logic;
        info_empty      : in     vl_logic;
        set_bus_error_irq: in     vl_logic;
        set_arbitration_lost_irq: in     vl_logic;
        arbitration_lost_capture: in     vl_logic_vector(4 downto 0);
        node_error_passive: in     vl_logic;
        node_error_active: in     vl_logic;
        rx_message_counter: in     vl_logic_vector(6 downto 0);
        reset_mode      : out    vl_logic;
        listen_only_mode: out    vl_logic;
        acceptance_filter_mode: out    vl_logic;
        self_test_mode  : out    vl_logic;
        clear_data_overrun: out    vl_logic;
        release_buffer  : out    vl_logic;
        abort_tx        : out    vl_logic;
        tx_request      : out    vl_logic;
        self_rx_request : out    vl_logic;
        single_shot_transmission: out    vl_logic;
        read_arbitration_lost_capture_reg: out    vl_logic;
        read_error_code_capture_reg: out    vl_logic;
        error_capture_code: in     vl_logic_vector(7 downto 0);
        baud_r_presc    : out    vl_logic_vector(5 downto 0);
        sync_jump_width : out    vl_logic_vector(1 downto 0);
        time_segment1   : out    vl_logic_vector(3 downto 0);
        time_segment2   : out    vl_logic_vector(2 downto 0);
        triple_sampling : out    vl_logic;
        error_warning_limit: out    vl_logic_vector(7 downto 0);
        we_rx_err_cnt   : out    vl_logic;
        we_tx_err_cnt   : out    vl_logic;
        extended_mode   : out    vl_logic;
        clkout          : out    vl_logic;
        acceptance_code_0: out    vl_logic_vector(7 downto 0);
        acceptance_mask_0: out    vl_logic_vector(7 downto 0);
        acceptance_code_1: out    vl_logic_vector(7 downto 0);
        acceptance_code_2: out    vl_logic_vector(7 downto 0);
        acceptance_code_3: out    vl_logic_vector(7 downto 0);
        acceptance_mask_1: out    vl_logic_vector(7 downto 0);
        acceptance_mask_2: out    vl_logic_vector(7 downto 0);
        acceptance_mask_3: out    vl_logic_vector(7 downto 0);
        tx_data_0       : out    vl_logic_vector(7 downto 0);
        tx_data_1       : out    vl_logic_vector(7 downto 0);
        tx_data_2       : out    vl_logic_vector(7 downto 0);
        tx_data_3       : out    vl_logic_vector(7 downto 0);
        tx_data_4       : out    vl_logic_vector(7 downto 0);
        tx_data_5       : out    vl_logic_vector(7 downto 0);
        tx_data_6       : out    vl_logic_vector(7 downto 0);
        tx_data_7       : out    vl_logic_vector(7 downto 0);
        tx_data_8       : out    vl_logic_vector(7 downto 0);
        tx_data_9       : out    vl_logic_vector(7 downto 0);
        tx_data_10      : out    vl_logic_vector(7 downto 0);
        tx_data_11      : out    vl_logic_vector(7 downto 0);
        tx_data_12      : out    vl_logic_vector(7 downto 0)
    );
end can_registers;
